
`include 'test_one.v'
`include 'test_three.v'
