module TEST_ONE(
  input rx,
  output tx
);

endmodule
